// Copyright (C) 2025  Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Altera and sold by Altera or its authorized distributors.  Please
// refer to the Altera Software License Subscription Agreements 
// on the Quartus Prime software download page.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 24.1std.0 Build 1077 03/04/2025 SC Lite Edition"
// CREATED		"Fri Sep 26 11:48:10 2025"

module seven_segment_decoder(
	D,
	S
);


input wire	[3:0] D;
output wire	[6:0] S;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;




assign	S[6] = D[3] | SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_2 & D[3];

assign	SYNTHESIZED_WIRE_80 = SYNTHESIZED_WIRE_81 & D[1];

assign	SYNTHESIZED_WIRE_79 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_83 =  ~D[3];

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_6 & D[2];

assign	SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_45 = SYNTHESIZED_WIRE_82 & SYNTHESIZED_WIRE_84;

assign	S[3] = SYNTHESIZED_WIRE_12 | SYNTHESIZED_WIRE_13;

assign	SYNTHESIZED_WIRE_18 = SYNTHESIZED_WIRE_83 | D[0];

assign	SYNTHESIZED_WIRE_76 = SYNTHESIZED_WIRE_15 & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_19 = D[3] | D[0];

assign	SYNTHESIZED_WIRE_75 = SYNTHESIZED_WIRE_17 & D[3];

assign	SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_18 & D[1];

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_19 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_31 = SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_22;

assign	S[5] = SYNTHESIZED_WIRE_23 | SYNTHESIZED_WIRE_24 | SYNTHESIZED_WIRE_25;

assign	SYNTHESIZED_WIRE_33 = SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_26 = SYNTHESIZED_WIRE_81 & D[1];

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_31 & SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_33 & D[2];

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_82 | D[2] | D[0];

assign	S[2] = SYNTHESIZED_WIRE_35 | SYNTHESIZED_WIRE_36 | SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_37 = SYNTHESIZED_WIRE_38 & SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_35 = D[0] & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_36 = SYNTHESIZED_WIRE_84 & D[3];

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_84 | SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_15 = D[1] | SYNTHESIZED_WIRE_45;

assign	SYNTHESIZED_WIRE_44 = D[0] & D[1];

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_52 = SYNTHESIZED_WIRE_48 & SYNTHESIZED_WIRE_83;

assign	S[1] = SYNTHESIZED_WIRE_50 | SYNTHESIZED_WIRE_51 | SYNTHESIZED_WIRE_52;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_81 & D[1];

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_55;

assign	SYNTHESIZED_WIRE_84 =  ~D[2];

assign	SYNTHESIZED_WIRE_50 = SYNTHESIZED_WIRE_56 & SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_82 =  ~D[1];

assign	SYNTHESIZED_WIRE_51 = D[0] & SYNTHESIZED_WIRE_82 & D[3];

assign	SYNTHESIZED_WIRE_81 =  ~D[0];

assign	SYNTHESIZED_WIRE_64 = SYNTHESIZED_WIRE_59 & SYNTHESIZED_WIRE_83;

assign	SYNTHESIZED_WIRE_17 = D[2] | D[1];

assign	SYNTHESIZED_WIRE_61 = D[0] & D[2];

assign	SYNTHESIZED_WIRE_59 = D[1] | SYNTHESIZED_WIRE_61;

assign	S[0] = SYNTHESIZED_WIRE_62 | SYNTHESIZED_WIRE_63 | SYNTHESIZED_WIRE_64;

assign	SYNTHESIZED_WIRE_66 = D[3] | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_66 & SYNTHESIZED_WIRE_82;

assign	SYNTHESIZED_WIRE_62 = SYNTHESIZED_WIRE_68 & SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_74 = SYNTHESIZED_WIRE_81 | SYNTHESIZED_WIRE_84;

assign	SYNTHESIZED_WIRE_73 = D[2] | SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_63 = SYNTHESIZED_WIRE_73 & D[1];

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_74 & D[1];

assign	S[4] = SYNTHESIZED_WIRE_75 | SYNTHESIZED_WIRE_76;

assign	SYNTHESIZED_WIRE_0 = SYNTHESIZED_WIRE_82 & D[2];

assign	SYNTHESIZED_WIRE_2 = SYNTHESIZED_WIRE_84 | D[1];

assign	SYNTHESIZED_WIRE_6 = SYNTHESIZED_WIRE_79 | SYNTHESIZED_WIRE_80;


endmodule
